module Hs(x,y,b,d);
input x,y;
output b,d;
assign s=x^y;
assign c = ~x&y;
endmodule